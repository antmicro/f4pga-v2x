(* blackbox *)
module GATE(
  input  wire I0,
  input  wire I1,
  output wire O
);

endmodule
